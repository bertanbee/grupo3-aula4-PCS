`include "mux_4x1_1bit.v"

module mux_4x1_16bit (
    input [15:0] I0, I1, I2, I3,
    input A0, A1,
    output [15:0] Q
);

    mux_4x1_1bit U0 (.I0(I0[0]), .I1(I1[0]), .I2(I2[0]), .I3(I3[0]), .A0(A0), .A1(A1), .Q(Q[0]));
    mux_4x1_1bit U1 (.I0(I0[1]), .I1(I1[1]), .I2(I2[1]), .I3(I3[1]), .A0(A0), .A1(A1), .Q(Q[1]));
    mux_4x1_1bit U2 (.I0(I0[2]), .I1(I1[2]), .I2(I2[2]), .I3(I3[2]), .A0(A0), .A1(A1), .Q(Q[2]));
    mux_4x1_1bit U3 (.I0(I0[3]), .I1(I1[3]), .I2(I2[3]), .I3(I3[3]), .A0(A0), .A1(A1), .Q(Q[3]));
    mux_4x1_1bit U4 (.I0(I0[4]), .I1(I1[4]), .I2(I2[4]), .I3(I3[4]), .A0(A0), .A1(A1), .Q(Q[4]));
    mux_4x1_1bit U5 (.I0(I0[5]), .I1(I1[5]), .I2(I2[5]), .I3(I3[5]), .A0(A0), .A1(A1), .Q(Q[5]));
    mux_4x1_1bit U6 (.I0(I0[6]), .I1(I1[6]), .I2(I2[6]), .I3(I3[6]), .A0(A0), .A1(A1), .Q(Q[6]));
    mux_4x1_1bit U7 (.I0(I0[7]), .I1(I1[7]), .I2(I2[7]), .I3(I3[7]), .A0(A0), .A1(A1), .Q(Q[7]));
    mux_4x1_1bit U8 (.I0(I0[8]), .I1(I1[8]), .I2(I2[8]), .I3(I3[8]), .A0(A0), .A1(A1), .Q(Q[8]));
    mux_4x1_1bit U9 (.I0(I0[9]), .I1(I1[9]), .I2(I2[9]), .I3(I3[9]), .A0(A0), .A1(A1), .Q(Q[9]));
    mux_4x1_1bit U10 (.I0(I0[10]), .I1(I1[10]), .I2(I2[10]), .I3(I3[10]), .A0(A0), .A1(A1), .Q(Q[10]));
    mux_4x1_1bit U11 (.I0(I0[11]), .I1(I1[11]), .I2(I2[11]), .I3(I3[11]), .A0(A0), .A1(A1), .Q(Q[11]));
    mux_4x1_1bit U12 (.I0(I0[12]), .I1(I1[12]), .I2(I2[12]), .I3(I3[12]), .A0(A0), .A1(A1), .Q(Q[12]));
    mux_4x1_1bit U13 (.I0(I0[13]), .I1(I1[13]), .I2(I2[13]), .I3(I3[13]), .A0(A0), .A1(A1), .Q(Q[13]));
    mux_4x1_1bit U14 (.I0(I0[14]), .I1(I1[14]), .I2(I2[14]), .I3(I3[14]), .A0(A0), .A1(A1), .Q(Q[14]));
    mux_4x1_1bit U15 (.I0(I0[15]), .I1(I1[15]), .I2(I2[15]), .I3(I3[15]), .A0(A0), .A1(A1), .Q(Q[15]));

endmodule